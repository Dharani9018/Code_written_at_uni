module sr_ff (
    input wire S,       // Set
    input wire R,       // Reset
    input wire clk,     // Clock
    input wire rst,     // Asynchronous reset
    output reg Q        // Output
);

    always @(posedge clk or posedge rst) begin
        if (rst)
            Q <= 1'b0;              // Async reset to 0
        else begin
            case ({S, R})
                2'b00: Q <= Q;      // No change
                2'b01: Q <= 1'b0;   // Reset
                2'b10: Q <= 1'b1;   // Set
                2'b11: Q <= 1'bx;   // Invalid (both high)
            endcase
        end
    end

endmodule

